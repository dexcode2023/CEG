LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY fullAdder1Bit IS 
	PORT
	(
		A :  IN  STD_LOGIC;
		B :  IN  STD_LOGIC;
		Ci :  IN  STD_LOGIC;
		S :  OUT  STD_LOGIC;
		Co :  OUT  STD_LOGIC
	);
END fullAdder1Bit;

ARCHITECTURE bdf_type OF fullAdder1Bit IS 

SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;


BEGIN 



SYNTHESIZED_WIRE_4 <= A XOR B;


S <= SYNTHESIZED_WIRE_4 XOR Ci;


Co <= SYNTHESIZED_WIRE_1 OR SYNTHESIZED_WIRE_2;


SYNTHESIZED_WIRE_2 <= Ci AND SYNTHESIZED_WIRE_4;


SYNTHESIZED_WIRE_1 <= A AND B;


END bdf_type;