
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY mux_8_2 IS
	PORT (
		a, b  : IN STD_LOGIC_VECTOR (7 downto 0);
		sel 		: IN STD_LOGIC;
		y 		: OUT STD_LOGIC_VECTOR (7 downto 0)
	);
END mux_8_2;

ARCHITECTURE struct OF mux_8_2 IS

COMPONENT mux_1_2 IS
	PORT (
		input : IN STD_LOGIC_VECTOR (1 downto 0);
		sel : IN STD_LOGIC;
		y : OUT STD_LOGIC
	);
END COMPONENT;

BEGIN

	MUX_0: mux_1_2
	PORT MAP (
		  input(0) => a(0),
		  input(1) => b(0),
		  sel => sel,
		  y => y(0) );

	MUX_1: mux_1_2
	PORT MAP (
		  input(0) => a(1),
		  input(1) => b(1),
		  sel => sel,
		  y => y(1) );

	MUX_2: mux_1_2
	PORT MAP (
		  input(0) => a(2),
		  input(1) => b(2),
		  sel => sel,
		  y => y(2) );

	MUX_3: mux_1_2
	PORT MAP (
		  input(0) => a(3),
		  input(1) => b(3),
		  sel => sel,
		  y => y(3) );

	MUX_4: mux_1_2
	PORT MAP (
		  input(0) => a(4),
		  input(1) => b(4),
		  sel => sel,
		  y => y(4) );

	MUX_5: mux_1_2
	PORT MAP (
		  input(0) => a(5),
		  input(1) => b(5),
		  sel => sel,
		  y => y(5) );
	
	MUX_6: mux_1_2
	PORT MAP (
		  input(0) => a(6),
		  input(1) => b(6),
		  sel => sel,
		  y => y(6) );

	MUX_7: mux_1_2
	PORT MAP (
		  input(0) => a(7),
		  input(1) => b(7),
		  sel => sel,
		  y => y(7) );

END struct;